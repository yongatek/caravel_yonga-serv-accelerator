magic
tech sky130A
magscale 1 2
timestamp 1635477528
<< nwell >>
rect 1066 357125 298854 357446
rect 1066 356037 298854 356603
rect 1066 354949 298854 355515
rect 1066 353861 298854 354427
rect 1066 352773 298854 353339
rect 1066 351685 298854 352251
rect 1066 350597 298854 351163
rect 1066 349509 298854 350075
rect 1066 348421 298854 348987
rect 1066 347333 298854 347899
rect 1066 346245 298854 346811
rect 1066 345157 298854 345723
rect 1066 344069 298854 344635
rect 1066 342981 298854 343547
rect 1066 341893 298854 342459
rect 1066 340805 298854 341371
rect 1066 339717 298854 340283
rect 1066 338629 298854 339195
rect 1066 337541 298854 338107
rect 1066 336453 298854 337019
rect 1066 335365 298854 335931
rect 1066 334277 298854 334843
rect 1066 333189 298854 333755
rect 1066 332101 298854 332667
rect 1066 331013 298854 331579
rect 1066 329925 298854 330491
rect 1066 328837 298854 329403
rect 1066 327749 298854 328315
rect 1066 326661 298854 327227
rect 1066 325573 298854 326139
rect 1066 324485 298854 325051
rect 1066 323397 298854 323963
rect 1066 322309 298854 322875
rect 1066 321221 298854 321787
rect 1066 320133 298854 320699
rect 1066 319045 298854 319611
rect 1066 317957 298854 318523
rect 1066 316869 298854 317435
rect 1066 315781 298854 316347
rect 1066 314693 298854 315259
rect 1066 313605 298854 314171
rect 1066 312517 298854 313083
rect 1066 311429 298854 311995
rect 1066 310341 298854 310907
rect 1066 309253 298854 309819
rect 1066 308165 298854 308731
rect 1066 307077 298854 307643
rect 1066 305989 298854 306555
rect 1066 304901 298854 305467
rect 1066 303813 298854 304379
rect 1066 302725 298854 303291
rect 1066 301637 298854 302203
rect 1066 300549 298854 301115
rect 1066 299461 298854 300027
rect 1066 298373 298854 298939
rect 1066 297285 298854 297851
rect 1066 296197 298854 296763
rect 1066 295109 298854 295675
rect 1066 294021 298854 294587
rect 1066 292933 298854 293499
rect 1066 291845 298854 292411
rect 1066 290757 298854 291323
rect 1066 289669 298854 290235
rect 1066 288581 298854 289147
rect 1066 287493 298854 288059
rect 1066 286405 298854 286971
rect 1066 285317 298854 285883
rect 1066 284229 298854 284795
rect 1066 283141 298854 283707
rect 1066 282053 298854 282619
rect 1066 280965 298854 281531
rect 1066 279877 298854 280443
rect 1066 278789 298854 279355
rect 1066 277701 298854 278267
rect 1066 276613 298854 277179
rect 1066 275525 298854 276091
rect 1066 274437 298854 275003
rect 1066 273349 298854 273915
rect 1066 272261 298854 272827
rect 1066 271173 298854 271739
rect 1066 270085 298854 270651
rect 1066 268997 298854 269563
rect 1066 267909 298854 268475
rect 1066 266821 298854 267387
rect 1066 265733 298854 266299
rect 1066 264645 298854 265211
rect 1066 263557 298854 264123
rect 1066 262469 298854 263035
rect 1066 261381 298854 261947
rect 1066 260293 298854 260859
rect 1066 259205 298854 259771
rect 1066 258117 298854 258683
rect 1066 257029 298854 257595
rect 1066 255941 298854 256507
rect 1066 254853 298854 255419
rect 1066 253765 298854 254331
rect 1066 252677 298854 253243
rect 1066 251589 298854 252155
rect 1066 250501 298854 251067
rect 1066 249413 298854 249979
rect 1066 248325 298854 248891
rect 1066 247237 298854 247803
rect 1066 246149 298854 246715
rect 1066 245061 298854 245627
rect 1066 243973 298854 244539
rect 1066 242885 298854 243451
rect 1066 241797 298854 242363
rect 1066 240709 298854 241275
rect 1066 239621 298854 240187
rect 1066 238533 298854 239099
rect 1066 237445 298854 238011
rect 1066 236357 298854 236923
rect 1066 235269 298854 235835
rect 1066 234181 298854 234747
rect 1066 233093 298854 233659
rect 1066 232005 298854 232571
rect 1066 230917 298854 231483
rect 1066 229829 298854 230395
rect 1066 228741 298854 229307
rect 1066 227653 298854 228219
rect 1066 226565 298854 227131
rect 1066 225477 298854 226043
rect 1066 224389 298854 224955
rect 1066 223301 298854 223867
rect 1066 222213 298854 222779
rect 1066 221125 298854 221691
rect 1066 220037 298854 220603
rect 1066 218949 298854 219515
rect 1066 217861 298854 218427
rect 1066 216773 298854 217339
rect 1066 215685 298854 216251
rect 1066 214597 298854 215163
rect 1066 213509 298854 214075
rect 1066 212421 298854 212987
rect 1066 211333 298854 211899
rect 1066 210245 298854 210811
rect 1066 209157 298854 209723
rect 1066 208069 298854 208635
rect 1066 206981 298854 207547
rect 1066 205893 298854 206459
rect 1066 204805 298854 205371
rect 1066 203717 298854 204283
rect 1066 202629 298854 203195
rect 1066 201541 298854 202107
rect 1066 200453 298854 201019
rect 1066 199365 298854 199931
rect 1066 198277 298854 198843
rect 1066 197189 298854 197755
rect 1066 196101 298854 196667
rect 1066 195013 298854 195579
rect 1066 193925 298854 194491
rect 1066 192837 298854 193403
rect 1066 191749 298854 192315
rect 1066 190661 298854 191227
rect 1066 189573 298854 190139
rect 1066 188485 298854 189051
rect 1066 187397 298854 187963
rect 1066 186309 298854 186875
rect 1066 185221 298854 185787
rect 1066 184133 298854 184699
rect 1066 183045 298854 183611
rect 1066 181957 298854 182523
rect 1066 180869 298854 181435
rect 1066 179781 298854 180347
rect 1066 178693 298854 179259
rect 1066 177605 298854 178171
rect 1066 176517 298854 177083
rect 1066 175429 298854 175995
rect 1066 174341 298854 174907
rect 1066 173253 298854 173819
rect 1066 172165 298854 172731
rect 1066 171077 298854 171643
rect 1066 169989 298854 170555
rect 1066 168901 298854 169467
rect 1066 167813 298854 168379
rect 1066 166725 298854 167291
rect 1066 165637 298854 166203
rect 1066 164549 298854 165115
rect 1066 163461 298854 164027
rect 1066 162373 298854 162939
rect 1066 161285 298854 161851
rect 1066 160197 298854 160763
rect 1066 159109 298854 159675
rect 1066 158021 298854 158587
rect 1066 156933 298854 157499
rect 1066 155845 298854 156411
rect 1066 154757 298854 155323
rect 1066 153669 298854 154235
rect 1066 152581 298854 153147
rect 1066 151493 298854 152059
rect 1066 150405 298854 150971
rect 1066 149317 298854 149883
rect 1066 148229 298854 148795
rect 1066 147141 298854 147707
rect 1066 146053 298854 146619
rect 1066 144965 298854 145531
rect 1066 143877 298854 144443
rect 1066 142789 298854 143355
rect 1066 141701 298854 142267
rect 1066 140613 298854 141179
rect 1066 139525 298854 140091
rect 1066 138437 298854 139003
rect 1066 137349 298854 137915
rect 1066 136261 298854 136827
rect 1066 135173 298854 135739
rect 1066 134085 298854 134651
rect 1066 132997 298854 133563
rect 1066 131909 298854 132475
rect 1066 130821 298854 131387
rect 1066 129733 298854 130299
rect 1066 128645 298854 129211
rect 1066 127557 298854 128123
rect 1066 126469 298854 127035
rect 1066 125381 298854 125947
rect 1066 124293 298854 124859
rect 1066 123205 298854 123771
rect 1066 122117 298854 122683
rect 1066 121029 298854 121595
rect 1066 119941 298854 120507
rect 1066 118853 298854 119419
rect 1066 117765 298854 118331
rect 1066 116677 298854 117243
rect 1066 115589 298854 116155
rect 1066 114501 298854 115067
rect 1066 113413 298854 113979
rect 1066 112325 298854 112891
rect 1066 111237 298854 111803
rect 1066 110149 298854 110715
rect 1066 109061 298854 109627
rect 1066 107973 298854 108539
rect 1066 106885 298854 107451
rect 1066 105797 298854 106363
rect 1066 104709 298854 105275
rect 1066 103621 298854 104187
rect 1066 102533 298854 103099
rect 1066 101445 298854 102011
rect 1066 100357 298854 100923
rect 1066 99269 298854 99835
rect 1066 98181 298854 98747
rect 1066 97093 298854 97659
rect 1066 96005 298854 96571
rect 1066 94917 298854 95483
rect 1066 93829 298854 94395
rect 1066 92741 298854 93307
rect 1066 91653 298854 92219
rect 1066 90565 298854 91131
rect 1066 89477 298854 90043
rect 1066 88389 298854 88955
rect 1066 87301 298854 87867
rect 1066 86213 298854 86779
rect 1066 85125 298854 85691
rect 1066 84037 298854 84603
rect 1066 82949 298854 83515
rect 1066 81861 298854 82427
rect 1066 80773 298854 81339
rect 1066 79685 298854 80251
rect 1066 78597 298854 79163
rect 1066 77509 298854 78075
rect 1066 76421 298854 76987
rect 1066 75333 298854 75899
rect 1066 74245 298854 74811
rect 1066 73157 298854 73723
rect 1066 72069 298854 72635
rect 1066 70981 298854 71547
rect 1066 69893 298854 70459
rect 1066 68805 298854 69371
rect 1066 67717 298854 68283
rect 1066 66629 298854 67195
rect 1066 65541 298854 66107
rect 1066 64453 298854 65019
rect 1066 63365 298854 63931
rect 1066 62277 298854 62843
rect 1066 61189 298854 61755
rect 1066 60101 298854 60667
rect 1066 59013 298854 59579
rect 1066 57925 298854 58491
rect 1066 56837 298854 57403
rect 1066 55749 298854 56315
rect 1066 54661 298854 55227
rect 1066 53573 298854 54139
rect 1066 52485 298854 53051
rect 1066 51397 298854 51963
rect 1066 50309 298854 50875
rect 1066 49221 298854 49787
rect 1066 48133 298854 48699
rect 1066 47045 298854 47611
rect 1066 45957 298854 46523
rect 1066 44869 298854 45435
rect 1066 43781 298854 44347
rect 1066 42693 298854 43259
rect 1066 41605 298854 42171
rect 1066 40517 298854 41083
rect 1066 39429 298854 39995
rect 1066 38341 298854 38907
rect 1066 37253 298854 37819
rect 1066 36165 298854 36731
rect 1066 35077 298854 35643
rect 1066 33989 298854 34555
rect 1066 32901 298854 33467
rect 1066 31813 298854 32379
rect 1066 30725 298854 31291
rect 1066 29637 298854 30203
rect 1066 28549 298854 29115
rect 1066 27461 298854 28027
rect 1066 26373 298854 26939
rect 1066 25285 298854 25851
rect 1066 24197 298854 24763
rect 1066 23109 298854 23675
rect 1066 22021 298854 22587
rect 1066 20933 298854 21499
rect 1066 19845 298854 20411
rect 1066 18757 298854 19323
rect 1066 17669 298854 18235
rect 1066 16581 298854 17147
rect 1066 15493 298854 16059
rect 1066 14405 298854 14971
rect 1066 13317 298854 13883
rect 1066 12229 298854 12795
rect 1066 11141 298854 11707
rect 1066 10053 298854 10619
rect 1066 8965 298854 9531
rect 1066 7877 298854 8443
rect 1066 6789 298854 7355
rect 1066 5701 298854 6267
rect 1066 4613 298854 5179
rect 1066 3525 298854 4091
rect 1066 2437 298854 3003
<< obsli1 >>
rect 1104 1377 298816 357425
<< obsm1 >>
rect 1104 756 298816 357456
<< metal2 >>
rect 1950 359200 2006 360000
rect 5814 359200 5870 360000
rect 9770 359200 9826 360000
rect 13726 359200 13782 360000
rect 17682 359200 17738 360000
rect 21638 359200 21694 360000
rect 25594 359200 25650 360000
rect 29550 359200 29606 360000
rect 33506 359200 33562 360000
rect 37462 359200 37518 360000
rect 41418 359200 41474 360000
rect 45282 359200 45338 360000
rect 49238 359200 49294 360000
rect 53194 359200 53250 360000
rect 57150 359200 57206 360000
rect 61106 359200 61162 360000
rect 65062 359200 65118 360000
rect 69018 359200 69074 360000
rect 72974 359200 73030 360000
rect 76930 359200 76986 360000
rect 80886 359200 80942 360000
rect 84842 359200 84898 360000
rect 88706 359200 88762 360000
rect 92662 359200 92718 360000
rect 96618 359200 96674 360000
rect 100574 359200 100630 360000
rect 104530 359200 104586 360000
rect 108486 359200 108542 360000
rect 112442 359200 112498 360000
rect 116398 359200 116454 360000
rect 120354 359200 120410 360000
rect 124310 359200 124366 360000
rect 128266 359200 128322 360000
rect 132130 359200 132186 360000
rect 136086 359200 136142 360000
rect 140042 359200 140098 360000
rect 143998 359200 144054 360000
rect 147954 359200 148010 360000
rect 151910 359200 151966 360000
rect 155866 359200 155922 360000
rect 159822 359200 159878 360000
rect 163778 359200 163834 360000
rect 167734 359200 167790 360000
rect 171690 359200 171746 360000
rect 175554 359200 175610 360000
rect 179510 359200 179566 360000
rect 183466 359200 183522 360000
rect 187422 359200 187478 360000
rect 191378 359200 191434 360000
rect 195334 359200 195390 360000
rect 199290 359200 199346 360000
rect 203246 359200 203302 360000
rect 207202 359200 207258 360000
rect 211158 359200 211214 360000
rect 215114 359200 215170 360000
rect 218978 359200 219034 360000
rect 222934 359200 222990 360000
rect 226890 359200 226946 360000
rect 230846 359200 230902 360000
rect 234802 359200 234858 360000
rect 238758 359200 238814 360000
rect 242714 359200 242770 360000
rect 246670 359200 246726 360000
rect 250626 359200 250682 360000
rect 254582 359200 254638 360000
rect 258538 359200 258594 360000
rect 262402 359200 262458 360000
rect 266358 359200 266414 360000
rect 270314 359200 270370 360000
rect 274270 359200 274326 360000
rect 278226 359200 278282 360000
rect 282182 359200 282238 360000
rect 286138 359200 286194 360000
rect 290094 359200 290150 360000
rect 294050 359200 294106 360000
rect 298006 359200 298062 360000
rect 1306 0 1362 800
rect 3974 0 4030 800
rect 6734 0 6790 800
rect 9402 0 9458 800
rect 12162 0 12218 800
rect 14922 0 14978 800
rect 17590 0 17646 800
rect 20350 0 20406 800
rect 23110 0 23166 800
rect 25778 0 25834 800
rect 28538 0 28594 800
rect 31298 0 31354 800
rect 33966 0 34022 800
rect 36726 0 36782 800
rect 39486 0 39542 800
rect 42154 0 42210 800
rect 44914 0 44970 800
rect 47582 0 47638 800
rect 50342 0 50398 800
rect 53102 0 53158 800
rect 55770 0 55826 800
rect 58530 0 58586 800
rect 61290 0 61346 800
rect 63958 0 64014 800
rect 66718 0 66774 800
rect 69478 0 69534 800
rect 72146 0 72202 800
rect 74906 0 74962 800
rect 77666 0 77722 800
rect 80334 0 80390 800
rect 83094 0 83150 800
rect 85854 0 85910 800
rect 88522 0 88578 800
rect 91282 0 91338 800
rect 93950 0 94006 800
rect 96710 0 96766 800
rect 99470 0 99526 800
rect 102138 0 102194 800
rect 104898 0 104954 800
rect 107658 0 107714 800
rect 110326 0 110382 800
rect 113086 0 113142 800
rect 115846 0 115902 800
rect 118514 0 118570 800
rect 121274 0 121330 800
rect 124034 0 124090 800
rect 126702 0 126758 800
rect 129462 0 129518 800
rect 132130 0 132186 800
rect 134890 0 134946 800
rect 137650 0 137706 800
rect 140318 0 140374 800
rect 143078 0 143134 800
rect 145838 0 145894 800
rect 148506 0 148562 800
rect 151266 0 151322 800
rect 154026 0 154082 800
rect 156694 0 156750 800
rect 159454 0 159510 800
rect 162214 0 162270 800
rect 164882 0 164938 800
rect 167642 0 167698 800
rect 170402 0 170458 800
rect 173070 0 173126 800
rect 175830 0 175886 800
rect 178498 0 178554 800
rect 181258 0 181314 800
rect 184018 0 184074 800
rect 186686 0 186742 800
rect 189446 0 189502 800
rect 192206 0 192262 800
rect 194874 0 194930 800
rect 197634 0 197690 800
rect 200394 0 200450 800
rect 203062 0 203118 800
rect 205822 0 205878 800
rect 208582 0 208638 800
rect 211250 0 211306 800
rect 214010 0 214066 800
rect 216678 0 216734 800
rect 219438 0 219494 800
rect 222198 0 222254 800
rect 224866 0 224922 800
rect 227626 0 227682 800
rect 230386 0 230442 800
rect 233054 0 233110 800
rect 235814 0 235870 800
rect 238574 0 238630 800
rect 241242 0 241298 800
rect 244002 0 244058 800
rect 246762 0 246818 800
rect 249430 0 249486 800
rect 252190 0 252246 800
rect 254950 0 255006 800
rect 257618 0 257674 800
rect 260378 0 260434 800
rect 263046 0 263102 800
rect 265806 0 265862 800
rect 268566 0 268622 800
rect 271234 0 271290 800
rect 273994 0 274050 800
rect 276754 0 276810 800
rect 279422 0 279478 800
rect 282182 0 282238 800
rect 284942 0 284998 800
rect 287610 0 287666 800
rect 290370 0 290426 800
rect 293130 0 293186 800
rect 295798 0 295854 800
rect 298558 0 298614 800
<< obsm2 >>
rect 1308 359144 1894 359258
rect 2062 359144 5758 359258
rect 5926 359144 9714 359258
rect 9882 359144 13670 359258
rect 13838 359144 17626 359258
rect 17794 359144 21582 359258
rect 21750 359144 25538 359258
rect 25706 359144 29494 359258
rect 29662 359144 33450 359258
rect 33618 359144 37406 359258
rect 37574 359144 41362 359258
rect 41530 359144 45226 359258
rect 45394 359144 49182 359258
rect 49350 359144 53138 359258
rect 53306 359144 57094 359258
rect 57262 359144 61050 359258
rect 61218 359144 65006 359258
rect 65174 359144 68962 359258
rect 69130 359144 72918 359258
rect 73086 359144 76874 359258
rect 77042 359144 80830 359258
rect 80998 359144 84786 359258
rect 84954 359144 88650 359258
rect 88818 359144 92606 359258
rect 92774 359144 96562 359258
rect 96730 359144 100518 359258
rect 100686 359144 104474 359258
rect 104642 359144 108430 359258
rect 108598 359144 112386 359258
rect 112554 359144 116342 359258
rect 116510 359144 120298 359258
rect 120466 359144 124254 359258
rect 124422 359144 128210 359258
rect 128378 359144 132074 359258
rect 132242 359144 136030 359258
rect 136198 359144 139986 359258
rect 140154 359144 143942 359258
rect 144110 359144 147898 359258
rect 148066 359144 151854 359258
rect 152022 359144 155810 359258
rect 155978 359144 159766 359258
rect 159934 359144 163722 359258
rect 163890 359144 167678 359258
rect 167846 359144 171634 359258
rect 171802 359144 175498 359258
rect 175666 359144 179454 359258
rect 179622 359144 183410 359258
rect 183578 359144 187366 359258
rect 187534 359144 191322 359258
rect 191490 359144 195278 359258
rect 195446 359144 199234 359258
rect 199402 359144 203190 359258
rect 203358 359144 207146 359258
rect 207314 359144 211102 359258
rect 211270 359144 215058 359258
rect 215226 359144 218922 359258
rect 219090 359144 222878 359258
rect 223046 359144 226834 359258
rect 227002 359144 230790 359258
rect 230958 359144 234746 359258
rect 234914 359144 238702 359258
rect 238870 359144 242658 359258
rect 242826 359144 246614 359258
rect 246782 359144 250570 359258
rect 250738 359144 254526 359258
rect 254694 359144 258482 359258
rect 258650 359144 262346 359258
rect 262514 359144 266302 359258
rect 266470 359144 270258 359258
rect 270426 359144 274214 359258
rect 274382 359144 278170 359258
rect 278338 359144 282126 359258
rect 282294 359144 286082 359258
rect 286250 359144 290038 359258
rect 290206 359144 293994 359258
rect 294162 359144 297950 359258
rect 298118 359144 298612 359258
rect 1308 856 298612 359144
rect 1418 734 3918 856
rect 4086 734 6678 856
rect 6846 734 9346 856
rect 9514 734 12106 856
rect 12274 734 14866 856
rect 15034 734 17534 856
rect 17702 734 20294 856
rect 20462 734 23054 856
rect 23222 734 25722 856
rect 25890 734 28482 856
rect 28650 734 31242 856
rect 31410 734 33910 856
rect 34078 734 36670 856
rect 36838 734 39430 856
rect 39598 734 42098 856
rect 42266 734 44858 856
rect 45026 734 47526 856
rect 47694 734 50286 856
rect 50454 734 53046 856
rect 53214 734 55714 856
rect 55882 734 58474 856
rect 58642 734 61234 856
rect 61402 734 63902 856
rect 64070 734 66662 856
rect 66830 734 69422 856
rect 69590 734 72090 856
rect 72258 734 74850 856
rect 75018 734 77610 856
rect 77778 734 80278 856
rect 80446 734 83038 856
rect 83206 734 85798 856
rect 85966 734 88466 856
rect 88634 734 91226 856
rect 91394 734 93894 856
rect 94062 734 96654 856
rect 96822 734 99414 856
rect 99582 734 102082 856
rect 102250 734 104842 856
rect 105010 734 107602 856
rect 107770 734 110270 856
rect 110438 734 113030 856
rect 113198 734 115790 856
rect 115958 734 118458 856
rect 118626 734 121218 856
rect 121386 734 123978 856
rect 124146 734 126646 856
rect 126814 734 129406 856
rect 129574 734 132074 856
rect 132242 734 134834 856
rect 135002 734 137594 856
rect 137762 734 140262 856
rect 140430 734 143022 856
rect 143190 734 145782 856
rect 145950 734 148450 856
rect 148618 734 151210 856
rect 151378 734 153970 856
rect 154138 734 156638 856
rect 156806 734 159398 856
rect 159566 734 162158 856
rect 162326 734 164826 856
rect 164994 734 167586 856
rect 167754 734 170346 856
rect 170514 734 173014 856
rect 173182 734 175774 856
rect 175942 734 178442 856
rect 178610 734 181202 856
rect 181370 734 183962 856
rect 184130 734 186630 856
rect 186798 734 189390 856
rect 189558 734 192150 856
rect 192318 734 194818 856
rect 194986 734 197578 856
rect 197746 734 200338 856
rect 200506 734 203006 856
rect 203174 734 205766 856
rect 205934 734 208526 856
rect 208694 734 211194 856
rect 211362 734 213954 856
rect 214122 734 216622 856
rect 216790 734 219382 856
rect 219550 734 222142 856
rect 222310 734 224810 856
rect 224978 734 227570 856
rect 227738 734 230330 856
rect 230498 734 232998 856
rect 233166 734 235758 856
rect 235926 734 238518 856
rect 238686 734 241186 856
rect 241354 734 243946 856
rect 244114 734 246706 856
rect 246874 734 249374 856
rect 249542 734 252134 856
rect 252302 734 254894 856
rect 255062 734 257562 856
rect 257730 734 260322 856
rect 260490 734 262990 856
rect 263158 734 265750 856
rect 265918 734 268510 856
rect 268678 734 271178 856
rect 271346 734 273938 856
rect 274106 734 276698 856
rect 276866 734 279366 856
rect 279534 734 282126 856
rect 282294 734 284886 856
rect 285054 734 287554 856
rect 287722 734 290314 856
rect 290482 734 293074 856
rect 293242 734 295742 856
rect 295910 734 298502 856
<< obsm3 >>
rect 4208 2143 297699 357441
<< metal4 >>
rect 4208 2128 4528 357456
rect 19568 2128 19888 357456
rect 34928 2128 35248 357456
rect 50288 2128 50608 357456
rect 65648 2128 65968 357456
rect 81008 2128 81328 357456
rect 96368 2128 96688 357456
rect 111728 2128 112048 357456
rect 127088 2128 127408 357456
rect 142448 2128 142768 357456
rect 157808 2128 158128 357456
rect 173168 2128 173488 357456
rect 188528 2128 188848 357456
rect 203888 2128 204208 357456
rect 219248 2128 219568 357456
rect 234608 2128 234928 357456
rect 249968 2128 250288 357456
rect 265328 2128 265648 357456
rect 280688 2128 281008 357456
rect 296048 2128 296368 357456
<< obsm4 >>
rect 24899 3571 34848 357101
rect 35328 3571 50208 357101
rect 50688 3571 65568 357101
rect 66048 3571 80928 357101
rect 81408 3571 96288 357101
rect 96768 3571 111648 357101
rect 112128 3571 127008 357101
rect 127488 3571 142368 357101
rect 142848 3571 157728 357101
rect 158208 3571 173088 357101
rect 173568 3571 188448 357101
rect 188928 3571 203808 357101
rect 204288 3571 219168 357101
rect 219648 3571 231965 357101
<< labels >>
rlabel metal2 s 1950 359200 2006 360000 6 io_oeb[0]
port 1 nsew signal output
rlabel metal2 s 80886 359200 80942 360000 6 io_oeb[10]
port 2 nsew signal output
rlabel metal2 s 88706 359200 88762 360000 6 io_oeb[11]
port 3 nsew signal output
rlabel metal2 s 96618 359200 96674 360000 6 io_oeb[12]
port 4 nsew signal output
rlabel metal2 s 104530 359200 104586 360000 6 io_oeb[13]
port 5 nsew signal output
rlabel metal2 s 112442 359200 112498 360000 6 io_oeb[14]
port 6 nsew signal output
rlabel metal2 s 120354 359200 120410 360000 6 io_oeb[15]
port 7 nsew signal output
rlabel metal2 s 128266 359200 128322 360000 6 io_oeb[16]
port 8 nsew signal output
rlabel metal2 s 136086 359200 136142 360000 6 io_oeb[17]
port 9 nsew signal output
rlabel metal2 s 143998 359200 144054 360000 6 io_oeb[18]
port 10 nsew signal output
rlabel metal2 s 151910 359200 151966 360000 6 io_oeb[19]
port 11 nsew signal output
rlabel metal2 s 9770 359200 9826 360000 6 io_oeb[1]
port 12 nsew signal output
rlabel metal2 s 159822 359200 159878 360000 6 io_oeb[20]
port 13 nsew signal output
rlabel metal2 s 167734 359200 167790 360000 6 io_oeb[21]
port 14 nsew signal output
rlabel metal2 s 175554 359200 175610 360000 6 io_oeb[22]
port 15 nsew signal output
rlabel metal2 s 183466 359200 183522 360000 6 io_oeb[23]
port 16 nsew signal output
rlabel metal2 s 191378 359200 191434 360000 6 io_oeb[24]
port 17 nsew signal output
rlabel metal2 s 199290 359200 199346 360000 6 io_oeb[25]
port 18 nsew signal output
rlabel metal2 s 207202 359200 207258 360000 6 io_oeb[26]
port 19 nsew signal output
rlabel metal2 s 215114 359200 215170 360000 6 io_oeb[27]
port 20 nsew signal output
rlabel metal2 s 222934 359200 222990 360000 6 io_oeb[28]
port 21 nsew signal output
rlabel metal2 s 230846 359200 230902 360000 6 io_oeb[29]
port 22 nsew signal output
rlabel metal2 s 17682 359200 17738 360000 6 io_oeb[2]
port 23 nsew signal output
rlabel metal2 s 238758 359200 238814 360000 6 io_oeb[30]
port 24 nsew signal output
rlabel metal2 s 246670 359200 246726 360000 6 io_oeb[31]
port 25 nsew signal output
rlabel metal2 s 254582 359200 254638 360000 6 io_oeb[32]
port 26 nsew signal output
rlabel metal2 s 262402 359200 262458 360000 6 io_oeb[33]
port 27 nsew signal output
rlabel metal2 s 270314 359200 270370 360000 6 io_oeb[34]
port 28 nsew signal output
rlabel metal2 s 278226 359200 278282 360000 6 io_oeb[35]
port 29 nsew signal output
rlabel metal2 s 286138 359200 286194 360000 6 io_oeb[36]
port 30 nsew signal output
rlabel metal2 s 294050 359200 294106 360000 6 io_oeb[37]
port 31 nsew signal output
rlabel metal2 s 25594 359200 25650 360000 6 io_oeb[3]
port 32 nsew signal output
rlabel metal2 s 33506 359200 33562 360000 6 io_oeb[4]
port 33 nsew signal output
rlabel metal2 s 41418 359200 41474 360000 6 io_oeb[5]
port 34 nsew signal output
rlabel metal2 s 49238 359200 49294 360000 6 io_oeb[6]
port 35 nsew signal output
rlabel metal2 s 57150 359200 57206 360000 6 io_oeb[7]
port 36 nsew signal output
rlabel metal2 s 65062 359200 65118 360000 6 io_oeb[8]
port 37 nsew signal output
rlabel metal2 s 72974 359200 73030 360000 6 io_oeb[9]
port 38 nsew signal output
rlabel metal2 s 5814 359200 5870 360000 6 io_out[0]
port 39 nsew signal output
rlabel metal2 s 84842 359200 84898 360000 6 io_out[10]
port 40 nsew signal output
rlabel metal2 s 92662 359200 92718 360000 6 io_out[11]
port 41 nsew signal output
rlabel metal2 s 100574 359200 100630 360000 6 io_out[12]
port 42 nsew signal output
rlabel metal2 s 108486 359200 108542 360000 6 io_out[13]
port 43 nsew signal output
rlabel metal2 s 116398 359200 116454 360000 6 io_out[14]
port 44 nsew signal output
rlabel metal2 s 124310 359200 124366 360000 6 io_out[15]
port 45 nsew signal output
rlabel metal2 s 132130 359200 132186 360000 6 io_out[16]
port 46 nsew signal output
rlabel metal2 s 140042 359200 140098 360000 6 io_out[17]
port 47 nsew signal output
rlabel metal2 s 147954 359200 148010 360000 6 io_out[18]
port 48 nsew signal output
rlabel metal2 s 155866 359200 155922 360000 6 io_out[19]
port 49 nsew signal output
rlabel metal2 s 13726 359200 13782 360000 6 io_out[1]
port 50 nsew signal output
rlabel metal2 s 163778 359200 163834 360000 6 io_out[20]
port 51 nsew signal output
rlabel metal2 s 171690 359200 171746 360000 6 io_out[21]
port 52 nsew signal output
rlabel metal2 s 179510 359200 179566 360000 6 io_out[22]
port 53 nsew signal output
rlabel metal2 s 187422 359200 187478 360000 6 io_out[23]
port 54 nsew signal output
rlabel metal2 s 195334 359200 195390 360000 6 io_out[24]
port 55 nsew signal output
rlabel metal2 s 203246 359200 203302 360000 6 io_out[25]
port 56 nsew signal output
rlabel metal2 s 211158 359200 211214 360000 6 io_out[26]
port 57 nsew signal output
rlabel metal2 s 218978 359200 219034 360000 6 io_out[27]
port 58 nsew signal output
rlabel metal2 s 226890 359200 226946 360000 6 io_out[28]
port 59 nsew signal output
rlabel metal2 s 234802 359200 234858 360000 6 io_out[29]
port 60 nsew signal output
rlabel metal2 s 21638 359200 21694 360000 6 io_out[2]
port 61 nsew signal output
rlabel metal2 s 242714 359200 242770 360000 6 io_out[30]
port 62 nsew signal output
rlabel metal2 s 250626 359200 250682 360000 6 io_out[31]
port 63 nsew signal output
rlabel metal2 s 258538 359200 258594 360000 6 io_out[32]
port 64 nsew signal output
rlabel metal2 s 266358 359200 266414 360000 6 io_out[33]
port 65 nsew signal output
rlabel metal2 s 274270 359200 274326 360000 6 io_out[34]
port 66 nsew signal output
rlabel metal2 s 282182 359200 282238 360000 6 io_out[35]
port 67 nsew signal output
rlabel metal2 s 290094 359200 290150 360000 6 io_out[36]
port 68 nsew signal output
rlabel metal2 s 298006 359200 298062 360000 6 io_out[37]
port 69 nsew signal output
rlabel metal2 s 29550 359200 29606 360000 6 io_out[3]
port 70 nsew signal output
rlabel metal2 s 37462 359200 37518 360000 6 io_out[4]
port 71 nsew signal output
rlabel metal2 s 45282 359200 45338 360000 6 io_out[5]
port 72 nsew signal output
rlabel metal2 s 53194 359200 53250 360000 6 io_out[6]
port 73 nsew signal output
rlabel metal2 s 61106 359200 61162 360000 6 io_out[7]
port 74 nsew signal output
rlabel metal2 s 69018 359200 69074 360000 6 io_out[8]
port 75 nsew signal output
rlabel metal2 s 76930 359200 76986 360000 6 io_out[9]
port 76 nsew signal output
rlabel metal2 s 293130 0 293186 800 6 irq[0]
port 77 nsew signal output
rlabel metal2 s 295798 0 295854 800 6 irq[1]
port 78 nsew signal output
rlabel metal2 s 298558 0 298614 800 6 irq[2]
port 79 nsew signal output
rlabel metal2 s 290370 0 290426 800 6 la_data_in
port 80 nsew signal input
rlabel metal4 s 4208 2128 4528 357456 6 vccd1
port 81 nsew power input
rlabel metal4 s 34928 2128 35248 357456 6 vccd1
port 81 nsew power input
rlabel metal4 s 65648 2128 65968 357456 6 vccd1
port 81 nsew power input
rlabel metal4 s 96368 2128 96688 357456 6 vccd1
port 81 nsew power input
rlabel metal4 s 127088 2128 127408 357456 6 vccd1
port 81 nsew power input
rlabel metal4 s 157808 2128 158128 357456 6 vccd1
port 81 nsew power input
rlabel metal4 s 188528 2128 188848 357456 6 vccd1
port 81 nsew power input
rlabel metal4 s 219248 2128 219568 357456 6 vccd1
port 81 nsew power input
rlabel metal4 s 249968 2128 250288 357456 6 vccd1
port 81 nsew power input
rlabel metal4 s 280688 2128 281008 357456 6 vccd1
port 81 nsew power input
rlabel metal4 s 19568 2128 19888 357456 6 vssd1
port 82 nsew ground input
rlabel metal4 s 50288 2128 50608 357456 6 vssd1
port 82 nsew ground input
rlabel metal4 s 81008 2128 81328 357456 6 vssd1
port 82 nsew ground input
rlabel metal4 s 111728 2128 112048 357456 6 vssd1
port 82 nsew ground input
rlabel metal4 s 142448 2128 142768 357456 6 vssd1
port 82 nsew ground input
rlabel metal4 s 173168 2128 173488 357456 6 vssd1
port 82 nsew ground input
rlabel metal4 s 203888 2128 204208 357456 6 vssd1
port 82 nsew ground input
rlabel metal4 s 234608 2128 234928 357456 6 vssd1
port 82 nsew ground input
rlabel metal4 s 265328 2128 265648 357456 6 vssd1
port 82 nsew ground input
rlabel metal4 s 296048 2128 296368 357456 6 vssd1
port 82 nsew ground input
rlabel metal2 s 1306 0 1362 800 6 wb_clk_i
port 83 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wb_rst_i
port 84 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_ack_o
port 85 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[0]
port 86 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 wbs_adr_i[10]
port 87 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 wbs_adr_i[11]
port 88 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 wbs_adr_i[12]
port 89 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 wbs_adr_i[13]
port 90 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 wbs_adr_i[14]
port 91 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 wbs_adr_i[15]
port 92 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 wbs_adr_i[16]
port 93 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 wbs_adr_i[17]
port 94 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 wbs_adr_i[18]
port 95 nsew signal input
rlabel metal2 s 184018 0 184074 800 6 wbs_adr_i[19]
port 96 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[1]
port 97 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 wbs_adr_i[20]
port 98 nsew signal input
rlabel metal2 s 200394 0 200450 800 6 wbs_adr_i[21]
port 99 nsew signal input
rlabel metal2 s 208582 0 208638 800 6 wbs_adr_i[22]
port 100 nsew signal input
rlabel metal2 s 216678 0 216734 800 6 wbs_adr_i[23]
port 101 nsew signal input
rlabel metal2 s 224866 0 224922 800 6 wbs_adr_i[24]
port 102 nsew signal input
rlabel metal2 s 233054 0 233110 800 6 wbs_adr_i[25]
port 103 nsew signal input
rlabel metal2 s 241242 0 241298 800 6 wbs_adr_i[26]
port 104 nsew signal input
rlabel metal2 s 249430 0 249486 800 6 wbs_adr_i[27]
port 105 nsew signal input
rlabel metal2 s 257618 0 257674 800 6 wbs_adr_i[28]
port 106 nsew signal input
rlabel metal2 s 265806 0 265862 800 6 wbs_adr_i[29]
port 107 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[2]
port 108 nsew signal input
rlabel metal2 s 273994 0 274050 800 6 wbs_adr_i[30]
port 109 nsew signal input
rlabel metal2 s 282182 0 282238 800 6 wbs_adr_i[31]
port 110 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_adr_i[3]
port 111 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 wbs_adr_i[4]
port 112 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 wbs_adr_i[5]
port 113 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 wbs_adr_i[6]
port 114 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 wbs_adr_i[7]
port 115 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 wbs_adr_i[8]
port 116 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 wbs_adr_i[9]
port 117 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_cyc_i
port 118 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[0]
port 119 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 wbs_dat_i[10]
port 120 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 wbs_dat_i[11]
port 121 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 wbs_dat_i[12]
port 122 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 wbs_dat_i[13]
port 123 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 wbs_dat_i[14]
port 124 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 wbs_dat_i[15]
port 125 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 wbs_dat_i[16]
port 126 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 wbs_dat_i[17]
port 127 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 wbs_dat_i[18]
port 128 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 wbs_dat_i[19]
port 129 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_i[1]
port 130 nsew signal input
rlabel metal2 s 194874 0 194930 800 6 wbs_dat_i[20]
port 131 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 wbs_dat_i[21]
port 132 nsew signal input
rlabel metal2 s 211250 0 211306 800 6 wbs_dat_i[22]
port 133 nsew signal input
rlabel metal2 s 219438 0 219494 800 6 wbs_dat_i[23]
port 134 nsew signal input
rlabel metal2 s 227626 0 227682 800 6 wbs_dat_i[24]
port 135 nsew signal input
rlabel metal2 s 235814 0 235870 800 6 wbs_dat_i[25]
port 136 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 wbs_dat_i[26]
port 137 nsew signal input
rlabel metal2 s 252190 0 252246 800 6 wbs_dat_i[27]
port 138 nsew signal input
rlabel metal2 s 260378 0 260434 800 6 wbs_dat_i[28]
port 139 nsew signal input
rlabel metal2 s 268566 0 268622 800 6 wbs_dat_i[29]
port 140 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_i[2]
port 141 nsew signal input
rlabel metal2 s 276754 0 276810 800 6 wbs_dat_i[30]
port 142 nsew signal input
rlabel metal2 s 284942 0 284998 800 6 wbs_dat_i[31]
port 143 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_i[3]
port 144 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 wbs_dat_i[4]
port 145 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_i[5]
port 146 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 wbs_dat_i[6]
port 147 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 wbs_dat_i[7]
port 148 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 wbs_dat_i[8]
port 149 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 wbs_dat_i[9]
port 150 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_o[0]
port 151 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 wbs_dat_o[10]
port 152 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 wbs_dat_o[11]
port 153 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 wbs_dat_o[12]
port 154 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 wbs_dat_o[13]
port 155 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 wbs_dat_o[14]
port 156 nsew signal output
rlabel metal2 s 156694 0 156750 800 6 wbs_dat_o[15]
port 157 nsew signal output
rlabel metal2 s 164882 0 164938 800 6 wbs_dat_o[16]
port 158 nsew signal output
rlabel metal2 s 173070 0 173126 800 6 wbs_dat_o[17]
port 159 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 wbs_dat_o[18]
port 160 nsew signal output
rlabel metal2 s 189446 0 189502 800 6 wbs_dat_o[19]
port 161 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_o[1]
port 162 nsew signal output
rlabel metal2 s 197634 0 197690 800 6 wbs_dat_o[20]
port 163 nsew signal output
rlabel metal2 s 205822 0 205878 800 6 wbs_dat_o[21]
port 164 nsew signal output
rlabel metal2 s 214010 0 214066 800 6 wbs_dat_o[22]
port 165 nsew signal output
rlabel metal2 s 222198 0 222254 800 6 wbs_dat_o[23]
port 166 nsew signal output
rlabel metal2 s 230386 0 230442 800 6 wbs_dat_o[24]
port 167 nsew signal output
rlabel metal2 s 238574 0 238630 800 6 wbs_dat_o[25]
port 168 nsew signal output
rlabel metal2 s 246762 0 246818 800 6 wbs_dat_o[26]
port 169 nsew signal output
rlabel metal2 s 254950 0 255006 800 6 wbs_dat_o[27]
port 170 nsew signal output
rlabel metal2 s 263046 0 263102 800 6 wbs_dat_o[28]
port 171 nsew signal output
rlabel metal2 s 271234 0 271290 800 6 wbs_dat_o[29]
port 172 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_o[2]
port 173 nsew signal output
rlabel metal2 s 279422 0 279478 800 6 wbs_dat_o[30]
port 174 nsew signal output
rlabel metal2 s 287610 0 287666 800 6 wbs_dat_o[31]
port 175 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 wbs_dat_o[3]
port 176 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 wbs_dat_o[4]
port 177 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 wbs_dat_o[5]
port 178 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 wbs_dat_o[6]
port 179 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 wbs_dat_o[7]
port 180 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 wbs_dat_o[8]
port 181 nsew signal output
rlabel metal2 s 107658 0 107714 800 6 wbs_dat_o[9]
port 182 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_sel_i[0]
port 183 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_sel_i[1]
port 184 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_sel_i[2]
port 185 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_sel_i[3]
port 186 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_stb_i
port 187 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_we_i
port 188 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 300000 360000
string LEFview TRUE
string GDS_FILE /project/openlane/subservient_wrapped/runs/subservient_wrapped/results/magic/subservient_wrapped.gds
string GDS_END 197621572
string GDS_START 865970
<< end >>

